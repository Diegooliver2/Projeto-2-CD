library ieee;
use ieee.std_logic_1164.all;

entity Processador is
port
	(
		SC : out std_logic_vector(10 downto 0)
	);
end Processador;